`timescale 1ns / 1ps

module test(
		input [2:0] a
    );


endmodule
